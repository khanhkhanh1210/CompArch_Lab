module lsu(
    input logic             i_clk,              // Clock
    input logic             i_rst,              // Reset

    input logic  [31:0]      i_lsu_addr,         // Address for data read/write
    input logic  [31:0]      i_st_data,          // Data to be stored
    input logic             i_lsu_wren,         // Write enable signal (1 if writing)

    output logic [31:0]     o_ld_data,          // Data read from memory
    output logic [31:0]     o_io_ledr,          // Output for red LEDs
    output logic [31:0]     o_io_ledg,          // Output for green LEDs

    output logic [6:0]      o_io_hex,           // Output for 7-segment displays
    output logic [31:0]     o_io_lcd,           // Output for the LCD register

    input logic  [31:0]      i_io_sw,            // Input for switches
    input logic  [3:0]       i_io_btn            // Input for buttons
);





endmodule