module decoder